library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sync is
	port (
		clk 				: in std_logic;
		reset				: in std_logic;
		vs_sig 			: out std_logic;
		hs_sig 			: out std_logic;
		pixel_data 	: out std_logic_vector(11 downto 0);
		pot : in std_logic_vector(11 downto 0)
	);
end entity sync;

architecture behavioral of sync is

	-- Note / R: bits 11:8 / G: bits 7:4 / B: bits 3:0 /  MSB:LSB ->
	constant red : std_logic_vector(11 downto 0) := X"F00";
	constant white : std_logic_vector(11 downto 0) := X"FFF";
	constant black : std_logic_vector(11 downto 0) := X"000";
	constant blue : std_logic_vector(11 downto 0) := X"00B";
	constant green : std_logic_vector(11 downto 0) := X"1A4";
	constant orange : std_logic_vector(11 downto 0) := X"F80";
	constant yellow : std_logic_vector(11 downto 0) := X"FD0";
	constant brown : std_logic_vector(11 downto 0) := X"643";
	
	type MY_MEM is array (0 to 72519) of std_logic_vector(11 downto 0);
	constant USA : MY_MEM := (X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"FFF", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B", X"00B");

	type vs_states is (V_FRONT_PORCH, V_SYNC, V_BACK_PORCH, DATA);
	signal current_vs_state, next_vs_state : vs_states;
	
	type hs_states is (H_FRONT_PORCH, H_SYNC, H_BACK_PORCH, P_DATA);
	signal current_hs_state, next_hs_state : hs_states;
	
	type my_horiz is range 0 to 799;
	
	signal x_pos : integer := 0;
	signal y_pos : integer := 0;
	signal next_x_pos : integer := 0;
	signal next_y_pos : integer := 0;
	signal count1 : integer := 0;
	signal count2 : integer := 0;
	signal count1_mod : integer := 0;
	signal count2_mod : integer := 0;
	signal m : std_logic := '0';
	signal pad_pos : integer := 0;
	signal pot_sig : integer := 0;
	
begin
	process(clk, reset, current_vs_state, count1, count2, current_hs_state, x_pos, y_pos) 
	begin
		if rising_edge(clk) then
			if reset = '0' then	
				current_vs_state <= V_FRONT_PORCH;
				current_hs_state <= H_FRONT_PORCH;
				count1 <= 0;
				count2 <= 0;
				x_pos <= 0;
				y_pos <= 0;
			else
				x_pos <= next_x_pos;
				y_pos <= next_y_pos;
				if m = '0' then
					count1 <= count1 + 1;
					count2 <= count2 + 1;
				else
					count1 <= 0;
					count2 <= 0;
				end if;
				current_vs_state <= next_vs_state;
				current_hs_state <= next_hs_state;
			end if;
		end if;
	end process;
	
	process(count1, current_vs_state, count1_mod)
	begin
		count1_mod <= count1 mod 420000;
		case current_vs_state is
			when V_FRONT_PORCH =>
				m <= '0';
				vs_sig <= '1';
				if count1_mod < 8000 then
					next_vs_state <= V_FRONT_PORCH;
				else
					next_vs_state <= V_SYNC;
				end if;
				
			when V_SYNC =>
				m <= '0';
				vs_sig <= '0';
				if count1_mod < 9600 then
					next_vs_state <= V_SYNC;
				else	
					next_vs_state <= V_BACK_PORCH;
				end if;
				
			when V_BACK_PORCH =>
				m <= '0';
				vs_sig <= '1';
				if count1_mod < 36000 then
					next_vs_state <= V_BACK_PORCH;
				else
					next_vs_state <= DATA;
				end if;
				
			when DATA =>
				vs_sig <= '1';
				if count1_mod < 420000 and count1_mod >= 36000 then
					next_vs_state <= DATA;
					m <= '0';
				else
					next_vs_state <= V_FRONT_PORCH;
					m <= '1';
				end if;
		end case;	
	end process;
	
	process(count2,count2_mod, x_pos, y_pos, current_hs_state, current_vs_state)
	begin
		count2_mod <= count2 mod 800;
		case current_hs_state is
			when H_FRONT_PORCH =>
				hs_sig <= '1';
				pixel_data <= black;
				next_x_pos <= 0;
				next_y_pos <= y_pos; 
				if count2_mod < 16 then
					next_hs_state <= H_FRONT_PORCH;
				else	
					next_hs_state <= H_SYNC;
				end if;
				
			when H_SYNC =>
				hs_sig <= '0';
				pixel_data <= black;
				next_x_pos <= 0;
				next_y_pos <= y_pos;
				if count2_mod < 112 then 
					next_hs_state <= H_SYNC;
				else	
					next_hs_state <= H_BACK_PORCH;
				end if;
				
			when H_BACK_PORCH =>
				hs_sig <= '1';
				pixel_data <= black;
				next_x_pos <= 0;
				if count2_mod < 160 then 
					next_hs_state <= H_BACK_PORCH;next_y_pos <= y_pos;
				else	
					next_hs_state <= P_DATA;
					next_y_pos <= y_pos + 1;
				end if;
				
			when P_DATA =>
				hs_sig <= '1';
				if count2_mod < 800 and count2_mod >= 160 then 
					next_hs_state <= P_DATA;
					next_y_pos <= y_pos;
					next_x_pos <= x_pos + 1;
				else	
					next_hs_state <= H_FRONT_PORCH;
					next_y_pos <= y_pos;
					next_x_pos <= x_pos;
				end if;
				if current_vs_state = V_FRONT_PORCH or current_vs_state = V_SYNC or current_vs_state = V_BACK_PORCH then
					pixel_data <= black;
					next_x_pos <= 0;
					next_y_pos <= 0;
				else
					next_y_pos <= y_pos;
					next_x_pos <= x_pos + 1;
				end if;	
				
				if y_pos < 480 and y_pos >474 then
					if x_pos >= pad_pos and x_pos < pad_pos + 40 then
						pixel_data <= brown;
					else
						pixel_data <= black;
					end if;
				else
					pixel_data <= black;
				end if;
				
		end case;
	end process;
	
	process(pot_sig) begin
		if(pot_sig > 3605) then
			pad_pos <= 600;
		else
			pad_pos <= pot_sig/6;
		end if;
	end process;
	
	pot_sig <= to_integer(unsigned(pot));
end architecture behavioral;